-------------------------------------------------------------------------------
-- Title      : TIE-50206, Exercise 08
-- Project    : 
-------------------------------------------------------------------------------
-- File       : adder.vhd
-- Author     : Jonas Nikula, Tuomas Huuki
-- Company    : TUT
-- Created    : 11.01.2016
-- Platform   : 
-- Standard   : VHDL'87
-------------------------------------------------------------------------------
-- Description: Controller for Wolfson WM8731 -audio codec
-------------------------------------------------------------------------------
-- Copyright (c) 2016 
-------------------------------------------------------------------------------
-- Revisions  :
-- Date         Version     Author          Description
-- 11.01.2016   1.0         nikulaj         Created
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity audio_ctrl is
    generic
    (
    );
    port
    (
    );
end audio_ctrl;

architecture rtl of audio_ctrl is
-- signal declarations go here
begin
-- logic goes here
end rtl;
