-------------------------------------------------------------------------------
-- Title      : TIE-50206, Exercise 09
-- Project    :
-------------------------------------------------------------------------------
-- File       : tb_audio_ctrl.vhd
-- Author     : Tuomas Huuki
-- Company    : TUT
-- Created    : 11.1.2016
-- Platform   :
-- Standard   : VHDL'93
-------------------------------------------------------------------------------
-- Description: Ninth excercise.
-------------------------------------------------------------------------------
-- Copyright (c) 2016
-------------------------------------------------------------------------------
-- Revisions  :
-- Date        Version  Author  Description
-- 11.1.2016   1.0      tuhu    Created
-------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity tb_audio_ctrl is
  generic(
    data_width_g    : integer := 16;
    step_w_r_g      : integer := 1;
    step_w_l_g      : integer := 4
  );
end tb_audio_ctrl;

architecture testbench of tb_audio_ctrl is
  
  component audio_ctrl is
    generic(
      ref_clk_freq_g  : integer := 18432000;
      sample_rate_g   : integer := 48000;
      data_width_g    : integer
    );
    
    port(
      clk             : in std_logic;
      rst_n           : in std_logic;
      left_data_in    : in std_logic_vector(data_width_g - 1 downto 0);
      right_data_in   : in std_logic_vector(data_width_g - 1 downto 0);
      aud_bclk_out    : out std_logic;
      aud_data_out    : out std_logic;
      aud_lrclk_out   : out std_logic
    );
  end component;
  
  component audio_codec_model is
  generic(
    data_width_g    : integer
  );
  port(
    rst_n           : in std_logic;
    aud_data_in     : in std_logic;
    aud_bclk_in     : in std_logic;
    aud_lrclk_in    : in std_logic;
    
    value_left_out  : out std_logic_vector(data_width_g - 1 downto 0);
    value_right_out : out std_logic_vector(data_width_g - 1 downto 0)
  );
  end component;

  component wave_gen is 
  generic (
    width_g             : integer;
    step_g              : integer := 1 
  );
  port(
    clk                 : in std_logic; 
    rst_n               : in std_logic; 
    sync_clear_in       : in std_logic; 
    value_out           : out std_logic_vector(width_g - 1 downto 0)
  );
  end component;
  
  constant clockrate_ns_c : time := 50 ns;
  
  signal clk              : std_logic := '0';
  signal rst_n            : std_logic := '0';
  signal sync_r           : std_logic := '0';
  signal left_data_in_r   : std_logic_vector(data_width_g - 1 downto 0);
  signal right_data_in_r  : std_logic_vector(data_width_g - 1 downto 0);
  signal aud_bclk_out_r   : std_logic;
  signal aud_data_out_r   : std_logic;
  signal aud_lrclk_out_r  : std_logic;
  signal left_data_out_r   : std_logic_vector(data_width_g - 1 downto 0);
  signal right_data_out_r  : std_logic_vector(data_width_g - 1 downto 0);
  
begin -- testbench
  i_acontrol : audio_ctrl
    generic map(
      data_width_g => data_width_g
    )
    port map(
      rst_n => rst_n,
      clk => clk,
      aud_data_out  => aud_data_out_r,
      aud_bclk_out  => aud_bclk_out_r,
      aud_lrclk_out => aud_lrclk_out_r,
      left_data_in => left_data_in_r,
      right_data_in => right_data_in_r    
    );
    
  i_amodel : audio_codec_model 
    generic map(
      data_width_g => data_width_g
    )
    port map(
      rst_n => rst_n,
      aud_data_in => aud_data_out_r,
      aud_bclk_in => aud_bclk_out_r,
      aud_lrclk_in => aud_lrclk_out_r,
      value_left_out => left_data_out_r,
      value_right_out => right_data_out_r
    );
  
  i_wavegen_left : wave_gen
    generic map(
      width_g => data_width_g,
      step_g => step_w_l_g
    )
    port map(
      clk => clk,
      rst_n => rst_n,
      sync_clear_in => sync_r,
      value_out => left_data_in_r
    ); 
    
  i_wavegen_right : wave_gen
    generic map(
      width_g => data_width_g,
      step_g => step_w_r_g
    )
    port map(
      clk => clk,
      rst_n => rst_n,
      sync_clear_in => sync_r,
      value_out => right_data_in_r
    ); 
    
  clk <= not clk after clockrate_ns_c/2; -- Create clock pulse.
  rst_n <= '1' after clockrate_ns_c * 4; -- Reset high after 4 pulses.
  
  data_generator : process(clk, rst_n)
  begin
    if(rst_n = '0') then
      -- Reset registers ..
    elsif(clk'event and clk = '1') then
      -- Generate data ..
    end if;
  end process data_generator;
  
end testbench;